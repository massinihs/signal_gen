module sine_lut #(
    parameter SAMPLES_PER_PERIOD = 200
)(  input  logic       clk,
    input  logic [7:0] index,
    output logic [11:0] value
);
	
    logic [11:0] arb_wave [0:SAMPLES_PER_PERIOD-1];

    // Read Logic (Synchronous Read)
    always @(posedge clk) begin
        value <= arb_wave[index];
    end

    // Array of signal
    initial begin
        arb_wave = '{
            // 0–49 noise
            12'd912, 12'd204, 12'd2253, 12'd2006, 12'd1828,
            12'd1143, 12'd839, 12'd712, 12'd3456, 12'd260,
            12'd244, 12'd767, 12'd1791, 12'd1905, 12'd217,
            12'd1628, 12'd3436, 12'd1805, 12'd3679, 12'd2278,
            12'd53,  12'd1307, 12'd3462, 12'd2787, 12'd2276,
            12'd1273, 12'd1763, 12'd2757, 12'd837,  12'd759,
            12'd3112, 12'd792,  12'd2940, 12'd2817, 12'd2166,
            12'd355,  12'd3763, 12'd1022, 12'd3100, 12'd645,
            12'd2401, 12'd2962, 12'd1575, 12'd569,  12'd375,
            12'd1866, 12'd2370, 12'd653,  12'd1907, 12'd827,

            // 50–99 high-frequency
            12'd2048, 12'd2664, 12'd2946, 12'd2741, 12'd2160,
            12'd1519, 12'd1164, 12'd1289, 12'd1825, 12'd2481,
            12'd2903, 12'd2862, 12'd2379, 12'd1717, 12'd1234,
            12'd1193, 12'd1615, 12'd2271, 12'd2807, 12'd2932,
            12'd2577, 12'd1936, 12'd1355, 12'd1150, 12'd1432,
            12'd2048, 12'd2664, 12'd2946, 12'd2741, 12'd2160,
            12'd1519, 12'd1164, 12'd1289, 12'd1825, 12'd2481,
            12'd2903, 12'd2862, 12'd2379, 12'd1717, 12'd1234,
            12'd1193, 12'd1615, 12'd2271, 12'd2807, 12'd2932,
            12'd2577, 12'd1936, 12'd1355, 12'd1150, 12'd1432,

            // 100–149 low-frequency
            12'd2048, 12'd2198, 12'd2346, 12'd2489, 12'd2626,
            12'd2753, 12'd2869, 12'd2972, 12'd3061, 12'd3133,
            12'd3189, 12'd3226, 12'd3245, 12'd3245, 12'd3226,
            12'd3189, 12'd3133, 12'd3061, 12'd2972, 12'd2869,
            12'd2753, 12'd2626, 12'd2489, 12'd2346, 12'd2198,
            12'd2048, 12'd1898, 12'd1750, 12'd1607, 12'd1470,
            12'd1343, 12'd1227, 12'd1124, 12'd1035, 12'd963,
            12'd907,  12'd870,  12'd851, 12'd851, 12'd870,
            12'd907,  12'd963, 12'd1035, 12'd1124, 12'd1227,
            12'd1343, 12'd1470, 12'd1607, 12'd1750, 12'd1898,

            // 150–199 medium-frequency
            12'd2048, 12'd2305, 12'd2527, 12'd2681, 12'd2746,
            12'd2713, 12'd2587, 12'd2385, 12'd2135, 12'd1874,
            12'd1637, 12'd1457, 12'd1361, 12'd1361, 12'd1457,
            12'd1637, 12'd1874, 12'd2135, 12'd2385, 12'd2587,
            12'd2713, 12'd2746, 12'd2681, 12'd2527, 12'd2305,
            12'd2048, 12'd1791, 12'd1569, 12'd1415, 12'd1350,
            12'd1383, 12'd1509, 12'd1711, 12'd1961, 12'd2222,
            12'd2459, 12'd2639, 12'd2735, 12'd2735, 12'd2639,
            12'd2459, 12'd2222, 12'd1961, 12'd1711, 12'd1509,
            12'd1383, 12'd1350, 12'd1415, 12'd1569, 12'd1791
        };
    end

endmodule
